module moduleName #(
    parameters
) (
    // BRANCH Flags
    output wire zero,
    output wire neg, // if in1 < in2, neg = 1, 0 otherwise
    output wire negu, // unsigned in1 and in2

);
    
endmodule