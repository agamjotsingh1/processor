module shift_left_1 (
	input wire [63:0] in,
	input wire in,

	output wire [63:0] out,
);
	
endmodule

module shift_left(
	input wire [63:0] in,
	input wire [63:0] amount, // shift amount
	output wire [63:0] out,
	output wire [63:0] medial, // intermediate results (used in multiplier)
);
	
endmodule
